** Profile: "SCHEMATIC1-OpAmpSim"  [ C:\Cadence\Hlektroniki3\opamp_hlek3\opamp_hlek3-pspicefiles\schematic1\opampsim.sim ] 

** Creating circuit file "OpAmpSim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../opamp_hlek3-pspicefiles/opamp_hlek3.lib" 
* From [PSPICE NETLIST] section of C:\SPB_DATA\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "C:\Cadence\SPB_17.2\tools\pspice\library\nomd.lib" 
.lib "C:\Cadence\SPB_17.2\tools\pspice\library\nom.lib" 

*Analysis directives: 
.AC DEC 40 1 1e+10
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
